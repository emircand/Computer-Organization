module concat (
    output [31:0] jump_pc,
    input [3:0] pc_plus_4,
    input [25:0] instruction
);
    or or1(jump_pc[31], pc_plus_4[3]);
    or or2(jump_pc[30], pc_plus_4[2]);
    or or3(jump_pc[29], pc_plus_4[1]);
    or or4(jump_pc[28], pc_plus_4[0]);
    or or5(jump_pc[27], instruction[25]);
    or or6(jump_pc[26], instruction[24]);
    or or7(jump_pc[25], instruction[23]);
    or or8(jump_pc[24], instruction[22]);
    or or9(jump_pc[23], instruction[21]);
    or or10(jump_pc[22], instruction[20]);
    or or11(jump_pc[21], instruction[19]);
    or or12(jump_pc[20], instruction[18]);
    or or13(jump_pc[19], instruction[17]);
    or or14(jump_pc[18], instruction[16]);
    or or15(jump_pc[17], instruction[15]);
    or or16(jump_pc[16], instruction[14]);
    or or17(jump_pc[15], instruction[13]);
    or or18(jump_pc[14], instruction[12]);
    or or19(jump_pc[13], instruction[11]);
    or or20(jump_pc[12], instruction[10]);
    or or21(jump_pc[11], instruction[9]);
    or or22(jump_pc[10], instruction[8]);
    or or23(jump_pc[9], instruction[7]);
    or or24(jump_pc[8], instruction[6]);
    or or25(jump_pc[7], instruction[5]);
    or or26(jump_pc[6], instruction[4]);
    or or27(jump_pc[5], instruction[3]);
    or or28(jump_pc[4], instruction[2]);
    or or29(jump_pc[3], instruction[1]);
    or or30(jump_pc[2], instruction[0]);
    or or31(jump_pc[1], 1'b0);
    or or32(jump_pc[0], 1'b0);
endmodule