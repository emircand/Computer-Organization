module not_32(
	output [31:0] res, 
	input [31:0] a
);

not not0 (res[0], a[0]);
not not1 (res[1], a[1]);
not not2 (res[2], a[2]);
not not3 (res[3], a[3]);
not not4 (res[4], a[4]);
not not5 (res[5], a[5]);
not not6 (res[6], a[6]);
not not7 (res[7], a[7]);
not not8 (res[8], a[8]);
not not9 (res[9], a[9]);
not not10 (res[10], a[10]);
not not11 (res[11], a[11]);
not not12 (res[12], a[12]);
not not13 (res[13], a[13]);
not not14 (res[14], a[14]);
not not15 (res[15], a[15]);
not not16 (res[16], a[16]);
not not17 (res[17], a[17]);
not not18 (res[18], a[18]);
not not19 (res[19], a[19]);
not not20 (res[20], a[20]);
not not21 (res[21], a[21]);
not not22 (res[22], a[22]);
not not23 (res[23], a[23]);
not not24 (res[24], a[24]);
not not25 (res[25], a[25]);
not not26 (res[26], a[26]);
not not27 (res[27], a[27]);
not not28 (res[28], a[28]);
not not29 (res[29], a[29]);
not not30 (res[30], a[30]);
not not31 (res[31], a[31]);

endmodule