module mux_6_6to1(input [2:0] s, input [5:0] d0, d1, d2, d3, d4, d5, output [5:0] y);
    mux_1_6to1 mux0(.s0(s[0]), .s1(s[1]), .s2(s[2]), .d0(d0[0]), .d1(d1[0]), .d2(d2[0]), .d3(d3[0]), .d4(d4[0]), .d5(d5[0]), .y(y[0]));
    mux_1_6to1 mux1(.s0(s[0]), .s1(s[1]), .s2(s[2]), .d0(d0[1]), .d1(d1[1]), .d2(d2[1]), .d3(d3[1]), .d4(d4[1]), .d5(d5[1]), .y(y[1]));
    mux_1_6to1 mux2(.s0(s[0]), .s1(s[1]), .s2(s[2]), .d0(d0[2]), .d1(d1[2]), .d2(d2[2]), .d3(d3[2]), .d4(d4[2]), .d5(d5[2]), .y(y[2]));
    mux_1_6to1 mux3(.s0(s[0]), .s1(s[1]), .s2(s[2]), .d0(d0[3]), .d1(d1[3]), .d2(d2[3]), .d3(d3[3]), .d4(d4[3]), .d5(d5[3]), .y(y[3]));
    mux_1_6to1 mux4(.s0(s[0]), .s1(s[1]), .s2(s[2]), .d0(d0[4]), .d1(d1[4]), .d2(d2[4]), .d3(d3[4]), .d4(d4[4]), .d5(d5[4]), .y(y[4]));
    mux_1_6to1 mux5(.s0(s[0]), .s1(s[1]), .s2(s[2]), .d0(d0[5]), .d1(d1[5]), .d2(d2[5]), .d3(d3[5]), .d4(d4[5]), .d5(d5[5]), .y(y[5]));
    mux_1_6to1 mux6(.s0(s[0]), .s1(s[1]), .s2(s[2]), .d0(d0[6]), .d1(d1[6]), .d2(d2[6]), .d3(d3[6]), .d4(d4[6]), .d5(d5[6]), .y(y[6]));
endmodule
